//==============================================================================
// Copyright (c) 2022 agithubber777
//------------------------------------------------------------------------------
// Module      : wm8731_top
// Description : WM8731 Control Top
// Author      : agithubber777
// Created     : 2022/05/31
//------------------------------------------------------------------------------
// Version Control Log:
//
// File$
// Revision$
// Author$
// Date$
//==============================================================================