//==============================================================================
// Copyright (c) 2022 agithubber777
//------------------------------------------------------------------------------
// Module      : wm8731_data
// Description : WM8731 Data Interface
// Author      : agithubber777
// Created     : 2022/05/31
//------------------------------------------------------------------------------
// Version Control Log:
//
// File$
// Revision$
// Author$
// Date$
//==============================================================================