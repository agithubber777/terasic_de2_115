//==============================================================================
// Copyright (C) 2023 agithubber777
//------------------------------------------------------------------------------
// File        : wm8731_top.sv
// Description : WM8731 Control Top
// Author      : agithubber777 (agit.hubber@gmail.com)
// Created     : 2023/02/17
//==============================================================================