//==============================================================================
// Copyright (c) 2022 agithubber777
//------------------------------------------------------------------------------
// Module      : wm8731_reg
// Description : WM8731 Config Register Control
// Author      : agithubber777
// Created     : 2022/05/31
//------------------------------------------------------------------------------
// Version Control Log:
//
// File$
// Revision$
// Author$
// Date$
//==============================================================================